library verilog;
use verilog.vl_types.all;
entity mips_pp_tb is
end mips_pp_tb;
