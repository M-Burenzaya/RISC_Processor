library verilog;
use verilog.vl_types.all;
entity slt2_tb is
    generic(
        clk_period      : integer := 10
    );
end slt2_tb;
