library verilog;
use verilog.vl_types.all;
entity registerfile32_tb is
    generic(
        clk_period      : integer := 10
    );
end registerfile32_tb;
