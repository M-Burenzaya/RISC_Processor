library verilog;
use verilog.vl_types.all;
entity signext_tb is
    generic(
        clk_period      : integer := 10
    );
end signext_tb;
