library verilog;
use verilog.vl_types.all;
entity mips_scp_tb is
end mips_scp_tb;
